library verilog;
use verilog.vl_types.all;
entity BeMicro_MAX10_top_vlg_check_tst is
    port(
        AD5681R_LDACn   : in     vl_logic;
        AD5681R_RSTn    : in     vl_logic;
        AD5681R_SCL     : in     vl_logic;
        AD5681R_SDA     : in     vl_logic;
        AD5681R_SYNCn   : in     vl_logic;
        ADT7420_SCL     : in     vl_logic;
        ADT7420_SDA     : in     vl_logic;
        ADXL362_CS      : in     vl_logic;
        ADXL362_MOSI    : in     vl_logic;
        ADXL362_SCLK    : in     vl_logic;
        EG_P1           : in     vl_logic;
        EG_P2           : in     vl_logic;
        EG_P3           : in     vl_logic;
        EG_P4           : in     vl_logic;
        EG_P5           : in     vl_logic;
        EG_P6           : in     vl_logic;
        EG_P7           : in     vl_logic;
        EG_P8           : in     vl_logic;
        EG_P9           : in     vl_logic;
        EG_P10          : in     vl_logic;
        EG_P11          : in     vl_logic;
        EG_P12          : in     vl_logic;
        EG_P13          : in     vl_logic;
        EG_P14          : in     vl_logic;
        EG_P15          : in     vl_logic;
        EG_P16          : in     vl_logic;
        EG_P17          : in     vl_logic;
        EG_P18          : in     vl_logic;
        EG_P19          : in     vl_logic;
        EG_P20          : in     vl_logic;
        EG_P21          : in     vl_logic;
        EG_P22          : in     vl_logic;
        EG_P23          : in     vl_logic;
        EG_P24          : in     vl_logic;
        EG_P25          : in     vl_logic;
        EG_P26          : in     vl_logic;
        EG_P27          : in     vl_logic;
        EG_P28          : in     vl_logic;
        EG_P29          : in     vl_logic;
        EG_P35          : in     vl_logic;
        EG_P36          : in     vl_logic;
        EG_P37          : in     vl_logic;
        EG_P38          : in     vl_logic;
        EG_P39          : in     vl_logic;
        EG_P40          : in     vl_logic;
        EG_P41          : in     vl_logic;
        EG_P42          : in     vl_logic;
        EG_P43          : in     vl_logic;
        EG_P44          : in     vl_logic;
        EG_P45          : in     vl_logic;
        EG_P46          : in     vl_logic;
        EG_P47          : in     vl_logic;
        EG_P48          : in     vl_logic;
        EG_P49          : in     vl_logic;
        EG_P50          : in     vl_logic;
        EG_P51          : in     vl_logic;
        EG_P52          : in     vl_logic;
        EG_P53          : in     vl_logic;
        EG_P54          : in     vl_logic;
        EG_P55          : in     vl_logic;
        EG_P56          : in     vl_logic;
        EG_P57          : in     vl_logic;
        EG_P58          : in     vl_logic;
        EG_P59          : in     vl_logic;
        EG_P60          : in     vl_logic;
        GPIO_01         : in     vl_logic;
        GPIO_02         : in     vl_logic;
        GPIO_03         : in     vl_logic;
        GPIO_04         : in     vl_logic;
        GPIO_05         : in     vl_logic;
        GPIO_06         : in     vl_logic;
        GPIO_07         : in     vl_logic;
        GPIO_08         : in     vl_logic;
        GPIO_09         : in     vl_logic;
        GPIO_10         : in     vl_logic;
        GPIO_11         : in     vl_logic;
        GPIO_12         : in     vl_logic;
        GPIO_A          : in     vl_logic;
        GPIO_B          : in     vl_logic;
        GPIO_J3_15      : in     vl_logic;
        GPIO_J3_16      : in     vl_logic;
        GPIO_J3_17      : in     vl_logic;
        GPIO_J3_18      : in     vl_logic;
        GPIO_J3_19      : in     vl_logic;
        GPIO_J3_20      : in     vl_logic;
        GPIO_J3_21      : in     vl_logic;
        GPIO_J3_22      : in     vl_logic;
        GPIO_J3_23      : in     vl_logic;
        GPIO_J3_24      : in     vl_logic;
        GPIO_J3_25      : in     vl_logic;
        GPIO_J3_26      : in     vl_logic;
        GPIO_J3_27      : in     vl_logic;
        GPIO_J3_28      : in     vl_logic;
        GPIO_J3_31      : in     vl_logic;
        GPIO_J3_32      : in     vl_logic;
        GPIO_J3_33      : in     vl_logic;
        GPIO_J3_34      : in     vl_logic;
        GPIO_J3_35      : in     vl_logic;
        GPIO_J3_36      : in     vl_logic;
        GPIO_J3_37      : in     vl_logic;
        GPIO_J3_38      : in     vl_logic;
        GPIO_J3_39      : in     vl_logic;
        GPIO_J3_40      : in     vl_logic;
        GPIO_J4_11      : in     vl_logic;
        GPIO_J4_12      : in     vl_logic;
        GPIO_J4_13      : in     vl_logic;
        GPIO_J4_14      : in     vl_logic;
        GPIO_J4_15      : in     vl_logic;
        GPIO_J4_16      : in     vl_logic;
        GPIO_J4_19      : in     vl_logic;
        GPIO_J4_20      : in     vl_logic;
        GPIO_J4_21      : in     vl_logic;
        GPIO_J4_22      : in     vl_logic;
        GPIO_J4_23      : in     vl_logic;
        GPIO_J4_24      : in     vl_logic;
        GPIO_J4_27      : in     vl_logic;
        GPIO_J4_28      : in     vl_logic;
        GPIO_J4_29      : in     vl_logic;
        GPIO_J4_30      : in     vl_logic;
        GPIO_J4_31      : in     vl_logic;
        GPIO_J4_32      : in     vl_logic;
        GPIO_J4_35      : in     vl_logic;
        GPIO_J4_36      : in     vl_logic;
        GPIO_J4_37      : in     vl_logic;
        GPIO_J4_38      : in     vl_logic;
        GPIO_J4_39      : in     vl_logic;
        GPIO_J4_40      : in     vl_logic;
        I2C_SCL         : in     vl_logic;
        I2C_SDA         : in     vl_logic;
        PMOD_A          : in     vl_logic_vector(3 downto 0);
        PMOD_B          : in     vl_logic_vector(3 downto 0);
        PMOD_C          : in     vl_logic_vector(3 downto 0);
        PMOD_D          : in     vl_logic_vector(3 downto 0);
        RESET_EXPn      : in     vl_logic;
        SDRAM_A         : in     vl_logic_vector(12 downto 0);
        SDRAM_BA        : in     vl_logic_vector(1 downto 0);
        SDRAM_CASn      : in     vl_logic;
        SDRAM_CKE       : in     vl_logic;
        SDRAM_CLK       : in     vl_logic;
        SDRAM_CSn       : in     vl_logic;
        SDRAM_DQ        : in     vl_logic_vector(15 downto 0);
        SDRAM_DQMH      : in     vl_logic;
        SDRAM_DQML      : in     vl_logic;
        SDRAM_RASn      : in     vl_logic;
        SDRAM_WEn       : in     vl_logic;
        SFLASH_DATA     : in     vl_logic;
        SFLASH_DCLK     : in     vl_logic;
        USER_LED        : in     vl_logic_vector(8 downto 1);
        sampler_rx      : in     vl_logic
    );
end BeMicro_MAX10_top_vlg_check_tst;
