library verilog;
use verilog.vl_types.all;
entity BeMicro_MAX10_top_vlg_vec_tst is
end BeMicro_MAX10_top_vlg_vec_tst;
