library verilog;
use verilog.vl_types.all;
entity BeMicro_MAX10_top is
    port(
        SYS_CLK         : in     vl_logic;
        USER_CLK        : in     vl_logic;
        AD5681R_LDACn   : out    vl_logic;
        AD5681R_RSTn    : out    vl_logic;
        AD5681R_SCL     : out    vl_logic;
        AD5681R_SDA     : out    vl_logic;
        AD5681R_SYNCn   : out    vl_logic;
        ADT7420_CT      : in     vl_logic;
        ADT7420_INT     : in     vl_logic;
        ADT7420_SCL     : inout  vl_logic;
        ADT7420_SDA     : inout  vl_logic;
        ADXL362_CS      : out    vl_logic;
        ADXL362_INT1    : in     vl_logic;
        ADXL362_INT2    : in     vl_logic;
        ADXL362_MISO    : in     vl_logic;
        ADXL362_MOSI    : out    vl_logic;
        ADXL362_SCLK    : out    vl_logic;
        SDRAM_A         : out    vl_logic_vector(12 downto 0);
        SDRAM_BA        : out    vl_logic_vector(1 downto 0);
        SDRAM_CASn      : out    vl_logic;
        SDRAM_CKE       : out    vl_logic;
        SDRAM_CLK       : out    vl_logic;
        SDRAM_CSn       : out    vl_logic;
        SDRAM_DQ        : inout  vl_logic_vector(15 downto 0);
        SDRAM_DQMH      : out    vl_logic;
        SDRAM_DQML      : out    vl_logic;
        SDRAM_RASn      : out    vl_logic;
        SDRAM_WEn       : out    vl_logic;
        SFLASH_ASDI     : in     vl_logic;
        SFLASH_CSn      : in     vl_logic;
        SFLASH_DATA     : inout  vl_logic;
        SFLASH_DCLK     : inout  vl_logic;
        AIN             : in     vl_logic_vector(7 downto 0);
        PB              : in     vl_logic_vector(4 downto 1);
        USER_LED        : out    vl_logic_vector(8 downto 1);
        EG_P1           : inout  vl_logic;
        EG_P10          : inout  vl_logic;
        EG_P11          : inout  vl_logic;
        EG_P12          : inout  vl_logic;
        EG_P13          : inout  vl_logic;
        EG_P14          : inout  vl_logic;
        EG_P15          : inout  vl_logic;
        EG_P16          : inout  vl_logic;
        EG_P17          : inout  vl_logic;
        EG_P18          : inout  vl_logic;
        EG_P19          : inout  vl_logic;
        EG_P2           : inout  vl_logic;
        EG_P20          : inout  vl_logic;
        EG_P21          : inout  vl_logic;
        EG_P22          : inout  vl_logic;
        EG_P23          : inout  vl_logic;
        EG_P24          : inout  vl_logic;
        EG_P25          : inout  vl_logic;
        EG_P26          : inout  vl_logic;
        EG_P27          : inout  vl_logic;
        EG_P28          : inout  vl_logic;
        EG_P29          : inout  vl_logic;
        EG_P3           : inout  vl_logic;
        EG_P35          : inout  vl_logic;
        EG_P36          : inout  vl_logic;
        EG_P37          : inout  vl_logic;
        EG_P38          : inout  vl_logic;
        EG_P39          : inout  vl_logic;
        EG_P4           : inout  vl_logic;
        EG_P40          : inout  vl_logic;
        EG_P41          : inout  vl_logic;
        EG_P42          : inout  vl_logic;
        EG_P43          : inout  vl_logic;
        EG_P44          : inout  vl_logic;
        EG_P45          : inout  vl_logic;
        EG_P46          : inout  vl_logic;
        EG_P47          : inout  vl_logic;
        EG_P48          : inout  vl_logic;
        EG_P49          : inout  vl_logic;
        EG_P5           : inout  vl_logic;
        EG_P50          : inout  vl_logic;
        EG_P51          : inout  vl_logic;
        EG_P52          : inout  vl_logic;
        EG_P53          : inout  vl_logic;
        EG_P54          : inout  vl_logic;
        EG_P55          : inout  vl_logic;
        EG_P56          : inout  vl_logic;
        EG_P57          : inout  vl_logic;
        EG_P58          : inout  vl_logic;
        EG_P59          : inout  vl_logic;
        EG_P6           : inout  vl_logic;
        EG_P60          : inout  vl_logic;
        EG_P7           : inout  vl_logic;
        EG_P8           : inout  vl_logic;
        EG_P9           : inout  vl_logic;
        EXP_PRESENT     : in     vl_logic;
        RESET_EXPn      : out    vl_logic;
        GPIO_01         : inout  vl_logic;
        GPIO_02         : inout  vl_logic;
        GPIO_03         : inout  vl_logic;
        GPIO_04         : inout  vl_logic;
        GPIO_05         : inout  vl_logic;
        GPIO_06         : inout  vl_logic;
        GPIO_07         : inout  vl_logic;
        GPIO_08         : inout  vl_logic;
        GPIO_09         : inout  vl_logic;
        GPIO_10         : inout  vl_logic;
        GPIO_11         : inout  vl_logic;
        GPIO_12         : inout  vl_logic;
        GPIO_A          : inout  vl_logic;
        GPIO_B          : inout  vl_logic;
        I2C_SCL         : inout  vl_logic;
        I2C_SDA         : inout  vl_logic;
        GPIO_J3_15      : inout  vl_logic;
        GPIO_J3_16      : inout  vl_logic;
        GPIO_J3_17      : inout  vl_logic;
        GPIO_J3_18      : inout  vl_logic;
        GPIO_J3_19      : inout  vl_logic;
        GPIO_J3_20      : inout  vl_logic;
        GPIO_J3_21      : inout  vl_logic;
        GPIO_J3_22      : inout  vl_logic;
        GPIO_J3_23      : inout  vl_logic;
        GPIO_J3_24      : inout  vl_logic;
        GPIO_J3_25      : inout  vl_logic;
        GPIO_J3_26      : inout  vl_logic;
        GPIO_J3_27      : inout  vl_logic;
        GPIO_J3_28      : inout  vl_logic;
        GPIO_J3_31      : inout  vl_logic;
        GPIO_J3_32      : inout  vl_logic;
        GPIO_J3_33      : inout  vl_logic;
        GPIO_J3_34      : inout  vl_logic;
        GPIO_J3_35      : inout  vl_logic;
        GPIO_J3_36      : inout  vl_logic;
        GPIO_J3_37      : inout  vl_logic;
        GPIO_J3_38      : inout  vl_logic;
        GPIO_J3_39      : inout  vl_logic;
        GPIO_J3_40      : inout  vl_logic;
        GPIO_J4_11      : inout  vl_logic;
        GPIO_J4_12      : inout  vl_logic;
        GPIO_J4_13      : inout  vl_logic;
        GPIO_J4_14      : inout  vl_logic;
        GPIO_J4_15      : inout  vl_logic;
        GPIO_J4_16      : inout  vl_logic;
        GPIO_J4_19      : inout  vl_logic;
        GPIO_J4_20      : inout  vl_logic;
        GPIO_J4_21      : inout  vl_logic;
        GPIO_J4_22      : inout  vl_logic;
        GPIO_J4_23      : inout  vl_logic;
        GPIO_J4_24      : inout  vl_logic;
        GPIO_J4_27      : inout  vl_logic;
        GPIO_J4_28      : inout  vl_logic;
        GPIO_J4_29      : inout  vl_logic;
        GPIO_J4_30      : inout  vl_logic;
        GPIO_J4_31      : inout  vl_logic;
        GPIO_J4_32      : inout  vl_logic;
        GPIO_J4_35      : inout  vl_logic;
        GPIO_J4_36      : inout  vl_logic;
        GPIO_J4_37      : inout  vl_logic;
        GPIO_J4_38      : inout  vl_logic;
        GPIO_J4_39      : inout  vl_logic;
        GPIO_J4_40      : inout  vl_logic;
        PMOD_A          : inout  vl_logic_vector(3 downto 0);
        PMOD_B          : inout  vl_logic_vector(3 downto 0);
        PMOD_C          : inout  vl_logic_vector(3 downto 0);
        PMOD_D          : inout  vl_logic_vector(3 downto 0)
    );
end BeMicro_MAX10_top;
